// Use UART_Rx to receive data from watch
// Store data in FIFO until special char is received
// Use UART_Tx to send FIFO data to esp32 until empty 


module WatchBase();

endmodule